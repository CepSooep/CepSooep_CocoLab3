module animationDraw (
  output reg oDone;
)