module fill
    (
        CLOCK_50,                       //  On Board 50 MHz
        // Your inputs and outputs here
        SW,
        KEY,                            // On Board Keys
        // The ports below are for the VGA output.  Do not change.
        VGA_CLK,                        //  VGA Clock
        VGA_HS,                         //  VGA H_SYNC
        VGA_VS,                         //  VGA V_SYNC
        VGA_BLANK_N,                        //  VGA BLANK
        VGA_SYNC_N,                     //  VGA SYNC
        VGA_R,                          //  VGA Red[9:0]
        VGA_G,                          //  VGA Green[9:0]
        VGA_B                           //  VGA Blue[9:0]
    );


    input           CLOCK_50;               //  50 MHz
    input   [3:0]   KEY;  
    input   [9:0] SW; //ixycoord,  icolor                 
    // Declare your inputs and outputs here
    // Do not change the following outputs
    output          VGA_CLK;                //  VGA Clock
    output          VGA_HS;                 //  VGA H_SYNC
    output          VGA_VS;                 //  VGA V_SYNC
    output          VGA_BLANK_N;                //  VGA BLANK
    output          VGA_SYNC_N;             //  VGA SYNC
    output  [7:0]   VGA_R;                  //  VGA Red[7:0] Changed from 10 to 8-bit DAC
    output  [7:0]   VGA_G;                  //  VGA Green[7:0]
    output  [7:0]   VGA_B;                  //  VGA Blue[7:0]
   
    wire resetn;
    assign resetn = KEY[0];
	wire [2:0] color;
    wire [7:0] x;
    wire [6:0] y;
	wire oPlot, oDone;
    wire writeEn; //iPlot
   
    part2 MAIN(.iResetn(resetn),
               .iPlotBox(writeEn),
               .iBlack(KEY[2]),
               .iColour(SW[9:7]),
               .iLoadX(KEY[3]),
               .iXY_Coord(KEY[1]),
               .iClock(CLOCK_50),
               .oX(x),
               .oY(y),
               .oColour(color),
               .oPlot(oPlot),
               .oDone(oDone));


    // Create the colour, x, y and writeEn wires that are inputs to the controller.
    
     // Create an Instance of a VGA controller - there can be only one!
    // Define the number of colours as well as the initial background
    // image file (.MIF) for the controller.
    vga_adapter VGA(
            .resetn(resetn),
            .clock(CLOCK_50),
            .colour(color),
            .x(x),
            .y(y),
            .plot(writeEn),
            /* Signals for the DAC to drive the monitor. */
            .VGA_R(VGA_R),
            .VGA_G(VGA_G),
            .VGA_B(VGA_B),
            .VGA_HS(VGA_HS),
            .VGA_VS(VGA_VS),
            .VGA_BLANK(VGA_BLANK_N),
            .VGA_SYNC(VGA_SYNC_N),
            .VGA_CLK(VGA_CLK));
        defparam VGA.RESOLUTION = "160x120";
        defparam VGA.MONOCHROME = "FALSE";
        defparam VGA.BITS_PER_COLOUR_CHANNEL = 1;
        defparam VGA.BACKGROUND_IMAGE = "black.mif";
           
    // Put your code here. Your code should produce signals x,y,colour and writeEn
    // for the VGA controller, in addition to any other functionality your design may require.
   
   
endmodule
